module ROM_128(
	input clk,
	input in_valid,
	input rst_n,
	output reg [23:0] w_r,
	output reg [23:0] w_i,
	output reg[1:0] state
);
////////////////////////////////////////////
// Internal signals
reg valid,next_valid;
reg [8:0] count,next_count;
////////////////////////////////////////////
// Next state logic
always @(*) begin
    if(in_valid || valid)next_count = count + 1;
    else next_count = count;
    
    if (count<9'd128) 
        state = 2'd0;
    else if (count >= 9'd128 && count < 9'd256)
        state = 2'd1;
    else if (count >= 9'd256 && count < 9'd384)
        state = 2'd2;
    else state = 2'd3;

	case(count)
	9'd256: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 000000000000000000000000;
	 next_valid = 1'b1;
	 end
	9'd257: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111111010;
	 next_valid = 1'b1;
	 end
	9'd258: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110011;
	 next_valid = 1'b1;
	 end
	9'd259: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111101101;
	 next_valid = 1'b1;
	 end
	9'd260: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111100111;
	 next_valid = 1'b1;
	 end
	9'd261: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111100001;
	 next_valid = 1'b1;
	 end
	9'd262: begin 
	 w_r = 24'b 000000000000000011111101;
	 w_i = 24'b 111111111111111111011010;
	 next_valid = 1'b1;
	 end
	9'd263: begin 
	 w_r = 24'b 000000000000000011111100;
	 w_i = 24'b 111111111111111111010100;
	 next_valid = 1'b1;
	 end
	9'd264: begin 
	 w_r = 24'b 000000000000000011111011;
	 w_i = 24'b 111111111111111111001110;
	 next_valid = 1'b1;
	 end
	9'd265: begin 
	 w_r = 24'b 000000000000000011111010;
	 w_i = 24'b 111111111111111111001000;
	 next_valid = 1'b1;
	 end
	9'd266: begin 
	 w_r = 24'b 000000000000000011111000;
	 w_i = 24'b 111111111111111111000010;
	 next_valid = 1'b1;
	 end
	9'd267: begin 
	 w_r = 24'b 000000000000000011110111;
	 w_i = 24'b 111111111111111110111100;
	 next_valid = 1'b1;
	 end
	9'd268: begin 
	 w_r = 24'b 000000000000000011110101;
	 w_i = 24'b 111111111111111110110110;
	 next_valid = 1'b1;
	 end
	9'd269: begin 
	 w_r = 24'b 000000000000000011110011;
	 w_i = 24'b 111111111111111110110000;
	 next_valid = 1'b1;
	 end
	9'd270: begin 
	 w_r = 24'b 000000000000000011110001;
	 w_i = 24'b 111111111111111110101010;
	 next_valid = 1'b1;
	 end
	9'd271: begin 
	 w_r = 24'b 000000000000000011101111;
	 w_i = 24'b 111111111111111110100100;
	 next_valid = 1'b1;
	 end
	9'd272: begin 
	 w_r = 24'b 000000000000000011101101;
	 w_i = 24'b 111111111111111110011110;
	 next_valid = 1'b1;
	 end
	9'd273: begin 
	 w_r = 24'b 000000000000000011101010;
	 w_i = 24'b 111111111111111110011000;
	 next_valid = 1'b1;
	 end
	9'd274: begin 
	 w_r = 24'b 000000000000000011100111;
	 w_i = 24'b 111111111111111110010011;
	 next_valid = 1'b1;
	 end
	9'd275: begin 
	 w_r = 24'b 000000000000000011100101;
	 w_i = 24'b 111111111111111110001101;
	 next_valid = 1'b1;
	 end
	9'd276: begin 
	 w_r = 24'b 000000000000000011100010;
	 w_i = 24'b 111111111111111110000111;
	 next_valid = 1'b1;
	 end
	9'd277: begin 
	 w_r = 24'b 000000000000000011011111;
	 w_i = 24'b 111111111111111110000010;
	 next_valid = 1'b1;
	 end
	9'd278: begin 
	 w_r = 24'b 000000000000000011011100;
	 w_i = 24'b 111111111111111101111100;
	 next_valid = 1'b1;
	 end
	9'd279: begin 
	 w_r = 24'b 000000000000000011011000;
	 w_i = 24'b 111111111111111101110111;
	 next_valid = 1'b1;
	 end
	9'd280: begin 
	 w_r = 24'b 000000000000000011010101;
	 w_i = 24'b 111111111111111101110010;
	 next_valid = 1'b1;
	 end
	9'd281: begin 
	 w_r = 24'b 000000000000000011010001;
	 w_i = 24'b 111111111111111101101101;
	 next_valid = 1'b1;
	 end
	9'd282: begin 
	 w_r = 24'b 000000000000000011001110;
	 w_i = 24'b 111111111111111101101000;
	 next_valid = 1'b1;
	 end
	9'd283: begin 
	 w_r = 24'b 000000000000000011001010;
	 w_i = 24'b 111111111111111101100011;
	 next_valid = 1'b1;
	 end
	9'd284: begin 
	 w_r = 24'b 000000000000000011000110;
	 w_i = 24'b 111111111111111101011110;
	 next_valid = 1'b1;
	 end
	9'd285: begin 
	 w_r = 24'b 000000000000000011000010;
	 w_i = 24'b 111111111111111101011001;
	 next_valid = 1'b1;
	 end
	9'd286: begin 
	 w_r = 24'b 000000000000000010111110;
	 w_i = 24'b 111111111111111101010100;
	 next_valid = 1'b1;
	 end
	9'd287: begin 
	 w_r = 24'b 000000000000000010111001;
	 w_i = 24'b 111111111111111101001111;
	 next_valid = 1'b1;
	 end
	9'd288: begin 
	 w_r = 24'b 000000000000000010110101;
	 w_i = 24'b 111111111111111101001011;
	 next_valid = 1'b1;
	 end
	9'd289: begin 
	 w_r = 24'b 000000000000000010110001;
	 w_i = 24'b 111111111111111101000111;
	 next_valid = 1'b1;
	 end
	9'd290: begin 
	 w_r = 24'b 000000000000000010101100;
	 w_i = 24'b 111111111111111101000010;
	 next_valid = 1'b1;
	 end
	9'd291: begin 
	 w_r = 24'b 000000000000000010100111;
	 w_i = 24'b 111111111111111100111110;
	 next_valid = 1'b1;
	 end
	9'd292: begin 
	 w_r = 24'b 000000000000000010100010;
	 w_i = 24'b 111111111111111100111010;
	 next_valid = 1'b1;
	 end
	9'd293: begin 
	 w_r = 24'b 000000000000000010011101;
	 w_i = 24'b 111111111111111100110110;
	 next_valid = 1'b1;
	 end
	9'd294: begin 
	 w_r = 24'b 000000000000000010011000;
	 w_i = 24'b 111111111111111100110010;
	 next_valid = 1'b1;
	 end
	9'd295: begin 
	 w_r = 24'b 000000000000000010010011;
	 w_i = 24'b 111111111111111100101111;
	 next_valid = 1'b1;
	 end
	9'd296: begin 
	 w_r = 24'b 000000000000000010001110;
	 w_i = 24'b 111111111111111100101011;
	 next_valid = 1'b1;
	 end
	9'd297: begin 
	 w_r = 24'b 000000000000000010001001;
	 w_i = 24'b 111111111111111100101000;
	 next_valid = 1'b1;
	 end
	9'd298: begin 
	 w_r = 24'b 000000000000000010000100;
	 w_i = 24'b 111111111111111100100100;
	 next_valid = 1'b1;
	 end
	9'd299: begin 
	 w_r = 24'b 000000000000000001111110;
	 w_i = 24'b 111111111111111100100001;
	 next_valid = 1'b1;
	 end
	9'd300: begin 
	 w_r = 24'b 000000000000000001111001;
	 w_i = 24'b 111111111111111100011110;
	 next_valid = 1'b1;
	 end
	9'd301: begin 
	 w_r = 24'b 000000000000000001110011;
	 w_i = 24'b 111111111111111100011011;
	 next_valid = 1'b1;
	 end
	9'd302: begin 
	 w_r = 24'b 000000000000000001101101;
	 w_i = 24'b 111111111111111100011001;
	 next_valid = 1'b1;
	 end
	9'd303: begin 
	 w_r = 24'b 000000000000000001101000;
	 w_i = 24'b 111111111111111100010110;
	 next_valid = 1'b1;
	 end
	9'd304: begin 
	 w_r = 24'b 000000000000000001100010;
	 w_i = 24'b 111111111111111100010011;
	 next_valid = 1'b1;
	 end
	9'd305: begin 
	 w_r = 24'b 000000000000000001011100;
	 w_i = 24'b 111111111111111100010001;
	 next_valid = 1'b1;
	 end
	9'd306: begin 
	 w_r = 24'b 000000000000000001010110;
	 w_i = 24'b 111111111111111100001111;
	 next_valid = 1'b1;
	 end
	9'd307: begin 
	 w_r = 24'b 000000000000000001010000;
	 w_i = 24'b 111111111111111100001101;
	 next_valid = 1'b1;
	 end
	9'd308: begin 
	 w_r = 24'b 000000000000000001001010;
	 w_i = 24'b 111111111111111100001011;
	 next_valid = 1'b1;
	 end
	9'd309: begin 
	 w_r = 24'b 000000000000000001000100;
	 w_i = 24'b 111111111111111100001001;
	 next_valid = 1'b1;
	 end
	9'd310: begin 
	 w_r = 24'b 000000000000000000111110;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	9'd311: begin 
	 w_r = 24'b 000000000000000000111000;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	9'd312: begin 
	 w_r = 24'b 000000000000000000110010;
	 w_i = 24'b 111111111111111100000101;
	 next_valid = 1'b1;
	 end
	9'd313: begin 
	 w_r = 24'b 000000000000000000101100;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	9'd314: begin 
	 w_r = 24'b 000000000000000000100110;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	9'd315: begin 
	 w_r = 24'b 000000000000000000011111;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	9'd316: begin 
	 w_r = 24'b 000000000000000000011001;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	9'd317: begin 
	 w_r = 24'b 000000000000000000010011;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	9'd318: begin 
	 w_r = 24'b 000000000000000000001101;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	9'd319: begin 
	 w_r = 24'b 000000000000000000000110;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	9'd320: begin 
	 w_r = 24'b 000000000000000000000000;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	9'd321: begin 
	 w_r = 24'b 111111111111111111111010;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	9'd322: begin 
	 w_r = 24'b 111111111111111111110011;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	9'd323: begin 
	 w_r = 24'b 111111111111111111101101;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	9'd324: begin 
	 w_r = 24'b 111111111111111111100111;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	9'd325: begin 
	 w_r = 24'b 111111111111111111100001;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	9'd326: begin 
	 w_r = 24'b 111111111111111111011010;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	9'd327: begin 
	 w_r = 24'b 111111111111111111010100;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	9'd328: begin 
	 w_r = 24'b 111111111111111111001110;
	 w_i = 24'b 111111111111111100000101;
	 next_valid = 1'b1;
	 end
	9'd329: begin 
	 w_r = 24'b 111111111111111111001000;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	9'd330: begin 
	 w_r = 24'b 111111111111111111000010;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	9'd331: begin 
	 w_r = 24'b 111111111111111110111100;
	 w_i = 24'b 111111111111111100001001;
	 next_valid = 1'b1;
	 end
	9'd332: begin 
	 w_r = 24'b 111111111111111110110110;
	 w_i = 24'b 111111111111111100001011;
	 next_valid = 1'b1;
	 end
	9'd333: begin 
	 w_r = 24'b 111111111111111110110000;
	 w_i = 24'b 111111111111111100001101;
	 next_valid = 1'b1;
	 end
	9'd334: begin 
	 w_r = 24'b 111111111111111110101010;
	 w_i = 24'b 111111111111111100001111;
	 next_valid = 1'b1;
	 end
	9'd335: begin 
	 w_r = 24'b 111111111111111110100100;
	 w_i = 24'b 111111111111111100010001;
	 next_valid = 1'b1;
	 end
	9'd336: begin 
	 w_r = 24'b 111111111111111110011110;
	 w_i = 24'b 111111111111111100010011;
	 next_valid = 1'b1;
	 end
	9'd337: begin 
	 w_r = 24'b 111111111111111110011000;
	 w_i = 24'b 111111111111111100010110;
	 next_valid = 1'b1;
	 end
	9'd338: begin 
	 w_r = 24'b 111111111111111110010011;
	 w_i = 24'b 111111111111111100011001;
	 next_valid = 1'b1;
	 end
	9'd339: begin 
	 w_r = 24'b 111111111111111110001101;
	 w_i = 24'b 111111111111111100011011;
	 next_valid = 1'b1;
	 end
	9'd340: begin 
	 w_r = 24'b 111111111111111110000111;
	 w_i = 24'b 111111111111111100011110;
	 next_valid = 1'b1;
	 end
	9'd341: begin 
	 w_r = 24'b 111111111111111110000010;
	 w_i = 24'b 111111111111111100100001;
	 next_valid = 1'b1;
	 end
	9'd342: begin 
	 w_r = 24'b 111111111111111101111100;
	 w_i = 24'b 111111111111111100100100;
	 next_valid = 1'b1;
	 end
	9'd343: begin 
	 w_r = 24'b 111111111111111101110111;
	 w_i = 24'b 111111111111111100101000;
	 next_valid = 1'b1;
	 end
	9'd344: begin 
	 w_r = 24'b 111111111111111101110010;
	 w_i = 24'b 111111111111111100101011;
	 next_valid = 1'b1;
	 end
	9'd345: begin 
	 w_r = 24'b 111111111111111101101101;
	 w_i = 24'b 111111111111111100101111;
	 next_valid = 1'b1;
	 end
	9'd346: begin 
	 w_r = 24'b 111111111111111101101000;
	 w_i = 24'b 111111111111111100110010;
	 next_valid = 1'b1;
	 end
	9'd347: begin 
	 w_r = 24'b 111111111111111101100011;
	 w_i = 24'b 111111111111111100110110;
	 next_valid = 1'b1;
	 end
	9'd348: begin 
	 w_r = 24'b 111111111111111101011110;
	 w_i = 24'b 111111111111111100111010;
	 next_valid = 1'b1;
	 end
	9'd349: begin 
	 w_r = 24'b 111111111111111101011001;
	 w_i = 24'b 111111111111111100111110;
	 next_valid = 1'b1;
	 end
	9'd350: begin 
	 w_r = 24'b 111111111111111101010100;
	 w_i = 24'b 111111111111111101000010;
	 next_valid = 1'b1;
	 end
	9'd351: begin 
	 w_r = 24'b 111111111111111101001111;
	 w_i = 24'b 111111111111111101000111;
	 next_valid = 1'b1;
	 end
	9'd352: begin 
	 w_r = 24'b 111111111111111101001011;
	 w_i = 24'b 111111111111111101001011;
	 next_valid = 1'b1;
	 end
	9'd353: begin 
	 w_r = 24'b 111111111111111101000111;
	 w_i = 24'b 111111111111111101001111;
	 next_valid = 1'b1;
	 end
	9'd354: begin 
	 w_r = 24'b 111111111111111101000010;
	 w_i = 24'b 111111111111111101010100;
	 next_valid = 1'b1;
	 end
	9'd355: begin 
	 w_r = 24'b 111111111111111100111110;
	 w_i = 24'b 111111111111111101011001;
	 next_valid = 1'b1;
	 end
	9'd356: begin 
	 w_r = 24'b 111111111111111100111010;
	 w_i = 24'b 111111111111111101011110;
	 next_valid = 1'b1;
	 end
	9'd357: begin 
	 w_r = 24'b 111111111111111100110110;
	 w_i = 24'b 111111111111111101100011;
	 next_valid = 1'b1;
	 end
	9'd358: begin 
	 w_r = 24'b 111111111111111100110010;
	 w_i = 24'b 111111111111111101101000;
	 next_valid = 1'b1;
	 end
	9'd359: begin 
	 w_r = 24'b 111111111111111100101111;
	 w_i = 24'b 111111111111111101101101;
	 next_valid = 1'b1;
	 end
	9'd360: begin 
	 w_r = 24'b 111111111111111100101011;
	 w_i = 24'b 111111111111111101110010;
	 next_valid = 1'b1;
	 end
	9'd361: begin 
	 w_r = 24'b 111111111111111100101000;
	 w_i = 24'b 111111111111111101110111;
	 next_valid = 1'b1;
	 end
	9'd362: begin 
	 w_r = 24'b 111111111111111100100100;
	 w_i = 24'b 111111111111111101111100;
	 next_valid = 1'b1;
	 end
	9'd363: begin 
	 w_r = 24'b 111111111111111100100001;
	 w_i = 24'b 111111111111111110000010;
	 next_valid = 1'b1;
	 end
	9'd364: begin 
	 w_r = 24'b 111111111111111100011110;
	 w_i = 24'b 111111111111111110000111;
	 next_valid = 1'b1;
	 end
	9'd365: begin 
	 w_r = 24'b 111111111111111100011011;
	 w_i = 24'b 111111111111111110001101;
	 next_valid = 1'b1;
	 end
	9'd366: begin 
	 w_r = 24'b 111111111111111100011001;
	 w_i = 24'b 111111111111111110010011;
	 next_valid = 1'b1;
	 end
	9'd367: begin 
	 w_r = 24'b 111111111111111100010110;
	 w_i = 24'b 111111111111111110011000;
	 next_valid = 1'b1;
	 end
	9'd368: begin 
	 w_r = 24'b 111111111111111100010011;
	 w_i = 24'b 111111111111111110011110;
	 next_valid = 1'b1;
	 end
	9'd369: begin 
	 w_r = 24'b 111111111111111100010001;
	 w_i = 24'b 111111111111111110100100;
	 next_valid = 1'b1;
	 end
	9'd370: begin 
	 w_r = 24'b 111111111111111100001111;
	 w_i = 24'b 111111111111111110101010;
	 next_valid = 1'b1;
	 end
	9'd371: begin 
	 w_r = 24'b 111111111111111100001101;
	 w_i = 24'b 111111111111111110110000;
	 next_valid = 1'b1;
	 end
	9'd372: begin 
	 w_r = 24'b 111111111111111100001011;
	 w_i = 24'b 111111111111111110110110;
	 next_valid = 1'b1;
	 end
	9'd373: begin 
	 w_r = 24'b 111111111111111100001001;
	 w_i = 24'b 111111111111111110111100;
	 next_valid = 1'b1;
	 end
	9'd374: begin 
	 w_r = 24'b 111111111111111100001000;
	 w_i = 24'b 111111111111111111000010;
	 next_valid = 1'b1;
	 end
	9'd375: begin 
	 w_r = 24'b 111111111111111100000110;
	 w_i = 24'b 111111111111111111001000;
	 next_valid = 1'b1;
	 end
	9'd376: begin 
	 w_r = 24'b 111111111111111100000101;
	 w_i = 24'b 111111111111111111001110;
	 next_valid = 1'b1;
	 end
	9'd377: begin 
	 w_r = 24'b 111111111111111100000100;
	 w_i = 24'b 111111111111111111010100;
	 next_valid = 1'b1;
	 end
	9'd378: begin 
	 w_r = 24'b 111111111111111100000011;
	 w_i = 24'b 111111111111111111011010;
	 next_valid = 1'b1;
	 end
	9'd379: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111100001;
	 next_valid = 1'b1;
	 end
	9'd380: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111100111;
	 next_valid = 1'b1;
	 end
	9'd381: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111101101;
	 next_valid = 1'b1;
	 end
	9'd382: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110011;
	 next_valid = 1'b1;
	 end
	9'd383: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111111010;
	 next_valid = 1'b0;
	 end
	default: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 000000000000000000000000;
	 next_valid = 1'b1;
	 end
	endcase
end
////////////////////////////////////////////
// State register
always@(posedge clk or negedge rst_n)begin
    if(~rst_n)begin
        count <= 0;
        valid <= 0;
    end
    else if(in_valid)
    begin
        count <= next_count;
        valid <= in_valid;
    end
    else if (valid)
    begin
        count <= next_count;
        valid <= next_valid;
    end
end
endmodule